// Reset signal interface.
// Used in ~reset_driver~ class.
interface reset_if(input logic clk);
    logic reset;
endinterface
