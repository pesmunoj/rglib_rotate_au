// Sequencer
// The sequencer is a mediator who establishes a connection between sequence and driver.

typedef uvm_sequencer#(reset_agent_seq_item_base)
    reset_agent_sequencer_base;
