typedef uvm_sequencer#(rglib_rotate_agent_seq_item)
    rglib_rotate_agent_sequencer;
