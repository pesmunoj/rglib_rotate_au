package reset_agent_pkg;

    import uvm_pkg::*;         // [UVM] package
    `include "uvm_macros.svh"  // [UVM] package

    `include "reset_agent_seq_item_base.sv"
    `include "reset_agent_sequence_base.sv"
    `include "reset_agent_sequencer_base.sv"
    `include "reset_agent_monitor_base.sv"
    `include "reset_agent_driver_base.sv"
    `include "reset_agent_base.sv"

endpackage
