
package rglib_rotate_tb_typedefs;
    import rglib_rotate_params_pkg::*;
    typedef logic [RGLIB_ROTATE_DATA_WIDTH-1:0]         rotate_data_t;
    typedef logic [RGLIB_ROTATE_ROTATE_STAGE_NUM-1:0]   rotate_val_t;
endpackage
